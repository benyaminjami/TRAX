module constants;
parameter T_empty = 3'bxxx;
parameter T_slash_down = 3'b001; 
parameter T_slash_up = 3'b010; 
parameter T_plus_vrt = 3'b011; 
parameter T_plus_hz = 3'b100;
parameter T_baskslash_up = 3'b101;
parameter T_backsalsh_down = 3'b110;
endmodule
