module TRAX(
	input 	rx,
	output	tx,
	input clock 
	);

parameter	b_height = 8'b01100100;
parameter	b_width = 8'b01100100;


parameter	s_IDLE = 4'b0000;
parameter	s_SET_Tile = 4'b0001;
parameter	s_SET_Board = 4'b0010;
parameter	s_WFIRST_Move = 4'b0011;
parameter	s_BFIRST_Move = 4'b0100;
parameter	s_SHIFT_Down = 4'b0101;
parameter 	s_SHIFT_Right = 4'b0110;
parameter	s_MANDATORY_Tile = 4'b0111;
parameter	s_FIND_Moves = 4'b1000;
parameter	s_SEND_Move = 4'b1001;

reg			set_color = 0;
reg			first_move = 0;
reg			r_color = 0;
reg [3:0]	r_SM_Main = 0;
reg [21:0] 	r_send_move;
reg			r_start_transmit;
reg			r_reset;
reg [21:0]	r_receive_move;
reg [2:0]	r_up_tile;
reg [2:0]	r_down_tile;
reg [2:0]	r_right_tile;
reg [2:0]	r_left_tile;
reg 		r_tile_check_start;
reg [5:0]	r_tile_type;
reg			r_R_Shift = 0;
reg			r_D_Shift = 0;
reg [21:0]	r_set_tile;
reg			r_mandatory_check = 0;
reg	[21:0] 	r_possible_moves[100:0];
integer		possible_moves_cnt = 0;
reg [2:0]	board[b_width:0][b_height:0];

integer		x_board = 2,y_board = 2;
integer		i,j;



wire [21:0] received_move;
tranceiver inst_tranceiver(
	.rx(rx),
	.move_in(r_send_move),
	.start_transmit(r_start_transmit),
	.clock(clock),
	.reset(r_reset),
	.tx(tx),
	.move_out(received_move),
	.end_receive(end_receive),
	.color(color)
	);
wire [5:0] tile_type;
tile_check inst_tile_check(
		.tile_type(tile_type),
		.endsignal(tile_check_end),
		.start_signal(r_tile_check_start),
		.up_tile(r_up_tile),
		.down_tile(r_down_tile),
		.right_tile(r_right_type),
		.left_tile(r_left_type),
		.clock()
		);

always @(posedge clock)
begin
	case(r_SM_Main)
	s_IDLE :
	begin
		r_start_transmit = 0;
		if(end_receive == 1)
		begin
			
			if(set_color == 0)
			begin
				r_color = color;
				set_color = 1;
				r_SM_Main = s_SET_Board;
				i = 0;
				j = 0;
			end
			else
			begin
				r_SM_Main = s_SET_Tile;
				r_set_tile = received_move;			
			end
		end
	end

	s_SET_Board:
	begin
		board[i][j] = 3'b000;
		i = i + 1;
		if(i == b_width)
		begin
			j = j + 1;
			i = 0;
		end
		if(j == b_height)
		begin
			if(r_color == 0)
				r_SM_Main = s_WFIRST_Move;
			else begin
				r_SM_Main = s_BFIRST_Move;
			end
		end
	end

	s_SET_Tile:
	begin
		if(tile_check_end == 1)
		begin
			r_tile_type = tile_type;
			if(received_move[21:20] == 1 && r_tile_type[4] == 1)
				board[ r_set_tile[19:10]] [r_set_tile[9:0]] = 3'b101;

			else if(r_set_tile[21:20] == 1 && r_tile_type[5] == 1)
				board[ r_set_tile[19:10]] [r_set_tile[9:0]] = 3'b110;

			else if(r_set_tile[21:20] == 0 && r_tile_type[0] == 1)
				board[ r_set_tile[19:10]] [r_set_tile[9:0]] = 3'b001;

			else if(r_set_tile[21:20] == 0 && r_tile_type[1] == 1)
				board[ r_set_tile[19:10]] [r_set_tile[9:0]] = 3'b010;

			else if(r_set_tile[21:20] == 2 && r_tile_type[2] == 1)
				board[ r_set_tile[19:10]] [r_set_tile[9:0]] = 3'b011;

			else if(r_set_tile[21:20] == 2 && r_tile_type[3] == 1)
				board[ r_set_tile[19:10]] [r_set_tile[9:0]] = 3'b100;

			if(r_set_tile[9:0] == 0)
				r_R_Shift = 1;
			if(r_set_tile[9:0] == x_board)
				x_board = x_board + 1;
			if(r_set_tile[19:10] == 0)
				r_D_Shift = 1;
			if(r_set_tile[19:10] == y_board)
				y_board = y_board + 1;
			r_SM_Main = s_SHIFT_Right;
			i = b_width - 1;
			j = 0;
			r_tile_check_start = 0;
		end
		r_down_tile = board[ r_set_tile[19:10] + 1] [r_set_tile[9:0]];
		r_right_tile = board[ r_set_tile[19:10]] [r_set_tile[9:0] + 1];
		if(r_set_tile[9:0] == 0)
			r_left_tile = 0;		
		else
			r_left_tile = board[ r_set_tile[19:10]] [r_set_tile[9:0] - 1];
		if(r_set_tile[19:10] == 0)
			r_up_tile = 0;
		else
			r_right_tile = board[ r_set_tile[19:10] - 1] [r_set_tile[9:0]];
		r_tile_check_start = 1;
	end

	s_WFIRST_Move:
	begin
		r_send_move = 3'b010;
		r_start_transmit = 1;
		r_SM_Main = s_IDLE;
	end

	s_BFIRST_Move:
	begin
		if(end_receive == 1)
		begin
			if(received_move[21:20] == 2)
				board[1][1] = 3'b011;
			else begin
				board[1][1] = 3'b010;
			end	
		end	
		r_SM_Main = s_FIND_Moves;
		i = 1;
		j = 0;
	end

	s_SHIFT_Right:
	begin
		if(r_R_Shift == 1)
		begin
			board[j][i] = board[j][i - 1];
			i = i - 1;
			if(i == 0)
			begin
				board[j][0] = 0;
				j = j + 1;
				i = b_width - 1;
			end
			if(j == b_height)
			begin
				r_R_Shift = 0;
			end
		end
		else begin
			j = b_height - 1;
			i = 0;
			r_SM_Main = s_SHIFT_Down;
		end
	end

	s_SHIFT_Down:
	begin
		if(r_D_Shift == 1)
		begin
			board[j][i] = board[j][i - 1];
			i = i - 1;
			if(i == 0)
			begin
				board[j][0] = 0;
				j = j + 1;
				i = b_height - 1;
			end
			if(j == b_width)
			begin
				r_D_Shift = 0;
			end
		end
		else begin
			r_SM_Main = s_MANDATORY_Tile;
			i = 0;
			j = 1;
		end
	end

	s_MANDATORY_Tile:
	begin
		if(tile_check_end == 1 && r_tile_check_start == 1)
		begin
			if(tile_type == 1)
			begin
				r_mandatory_check = 1;
				board[i][j] = 1;
			end
			if(tile_type == 2)
			begin
				r_mandatory_check = 1;
				board[i][j] = 2;
			end
			if(tile_type == 4)
			begin
				r_mandatory_check = 1;
				board[i][j] = 3;
			end
			if(tile_type == 8)
			begin
				r_mandatory_check = 1;
				board[i][j] = 4;
			end
			if(tile_type == 16)
			begin
				r_mandatory_check = 1;
				board[i][j] = 5;
			end
			if(tile_type == 32)
			begin
				r_mandatory_check = 1;
				board[i][j] = 6;
			end			
			r_tile_check_start = 0;
			j = j + 1;
			if(j == b_width)
			begin
				j = 0;
				i = i + 1;
			end
			if(i == b_height)
			begin
				if(r_mandatory_check == 1)
				begin
					i = 0;
					j = 1;
					r_mandatory_check = 0;
				end
				else begin
					i = 1;
					j = 0;
					r_SM_Main = s_FIND_Moves;
				end
			end
		end
		r_down_tile = board[i + 1] [j];
		r_right_tile = board[i] [j + 1];
		if(j == 0)
			r_left_tile = 0;		
		else
			r_left_tile = board[i] [j - 1];
		if(i == 0)
			r_up_tile = 0;
		else
			r_right_tile = board[i - 1] [j];
		if(board[i][j] != 0)
		begin
			j = j + 1;
			if(j == b_width)
			begin
				j = 0;
				i = i + 1;
			end
		end
		else
			r_tile_check_start = 1;
	end

	s_FIND_Moves:
	begin
		if(tile_check_end == 1 && r_tile_check_start == 1)
		begin
			if(tile_type[0] == 1)
			begin
				r_possible_moves[possible_moves_cnt][9:0] = j;
				r_possible_moves[possible_moves_cnt][19:10] = i;
				r_possible_moves[possible_moves_cnt][21:20] = 0;
				possible_moves_cnt = possible_moves_cnt + 1;
			end
			if(tile_type[1] == 1)
			begin
				r_possible_moves[possible_moves_cnt][9:0] = j;
				r_possible_moves[possible_moves_cnt][19:10] = i;
				r_possible_moves[possible_moves_cnt][21:20] = 0;
				possible_moves_cnt = possible_moves_cnt + 1;
			end
			if(tile_type[2] == 1)
			begin
				r_possible_moves[possible_moves_cnt][9:0] = j;
				r_possible_moves[possible_moves_cnt][19:10] = i;
				r_possible_moves[possible_moves_cnt][21:20] = 1;
				possible_moves_cnt = possible_moves_cnt + 1;
			end
			if(tile_type[3] == 1)
			begin
				r_possible_moves[possible_moves_cnt][9:0] = j;
				r_possible_moves[possible_moves_cnt][19:10] = i;
				r_possible_moves[possible_moves_cnt][21:20] = 1;
				possible_moves_cnt = possible_moves_cnt + 1;
			end
			if(tile_type[4] == 1)
			begin
				r_possible_moves[possible_moves_cnt][9:0] = j;
				r_possible_moves[possible_moves_cnt][19:10] = i;
				r_possible_moves[possible_moves_cnt][21:20] = 2;
				possible_moves_cnt = possible_moves_cnt + 1;
			end
			if(tile_type[5] == 1)
			begin
				r_possible_moves[possible_moves_cnt][9:0] = j;
				r_possible_moves[possible_moves_cnt][19:10] = i;
				r_possible_moves[possible_moves_cnt][21:20] = 2;
				possible_moves_cnt = possible_moves_cnt + 1;
			end			
			r_tile_check_start = 0;
			j = j + 1;
			if(j == b_width)
			begin
				j = 0;
				i = i + 1;
			end
			if(i == b_height)
			begin
				r_SM_Main = s_SEND_Move;
			end
		end
		r_down_tile = board[i + 1] [j];
		r_right_tile = board[i] [j + 1];
		if(j == 0)
			r_left_tile = 0;		
		else
			r_left_tile = board[i] [j - 1];
		if(i == 0)
			r_up_tile = 0;
		else
			r_right_tile = board[i - 1] [j];
		if(board[i][j] != 0)
		begin
			j = j + 1;
			if(j == b_width)
			begin
				j = 0;
				i = i + 1;
			end
		end
		else
			r_tile_check_start = 1;
	end

	s_SEND_Move:
	begin
		r_send_move = r_possible_moves[0];
		r_start_transmit = 1;
		possible_moves_cnt = 0;
		r_SM_Main = s_IDLE;
	end

	default
		r_SM_Main = s_IDLE;

	endcase
end
endmodule
