module find_moves(
		output	[2099:0]	moves,
		output			end_signal,
		input			start_signal,
		input	[29999:0]	board,
		input			clock
		}

endmodule
