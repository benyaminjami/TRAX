module TRAX;

endmodule
