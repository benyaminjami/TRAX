module board_shift(
		output	[29999:0]	shifted_board,
		output			end_signal,
		input	[29999:0]	board,
		input			start_signal,
		input			right_shift,
		input			down_shift,
		input 			clock
		);

endmodule
