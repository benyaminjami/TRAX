module tile_check(
		output	[5:0]	tile_type,
		output		end_signal,
		input		start_signal,
		input	[2:0]	up_tile,
		input	[2:0]	down_tile,
		input	[2:0]	right_tile,
		input	[2:0]	left_tile
		);

endmodule
